
module issp_char (
	source);	

	output	[7:0]	source;
endmodule
