
module issp_position (
	source);	

	output	[6:0]	source;
endmodule
